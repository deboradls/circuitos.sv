module codprior3x8 (
    port_list
);
    
endmodule